magic
tech scmos
timestamp 1644280066
<< nwell >>
rect -5 -1 56 33
<< polysilicon >>
rect 5 24 7 26
rect 15 24 17 26
rect 24 24 26 26
rect 44 24 46 26
rect 5 -39 7 0
rect 15 -39 17 0
rect 24 -39 26 0
rect 44 -39 46 0
rect 5 -45 7 -43
rect 15 -45 17 -43
rect 24 -45 26 -43
rect 44 -45 46 -43
<< ndiffusion >>
rect 4 -43 5 -39
rect 7 -43 15 -39
rect 17 -43 24 -39
rect 26 -43 27 -39
rect 43 -43 44 -39
rect 46 -43 47 -39
<< pdiffusion >>
rect 4 0 5 24
rect 7 0 9 24
rect 13 0 15 24
rect 17 0 19 24
rect 23 0 24 24
rect 26 0 27 24
rect 43 0 44 24
rect 46 0 47 24
<< metal1 >>
rect -1 28 3 32
rect 7 28 11 32
rect 15 28 19 32
rect 23 28 27 32
rect 31 28 35 32
rect 9 24 13 28
rect 27 24 31 28
rect 39 24 43 32
rect 47 28 52 32
rect 0 -3 4 0
rect 19 -3 23 0
rect 0 -7 34 -3
rect -5 -14 1 -10
rect 30 -18 34 -7
rect 47 -18 51 0
rect -5 -22 11 -18
rect 30 -22 40 -18
rect 47 -22 56 -18
rect -5 -30 20 -26
rect 30 -27 34 -22
rect 27 -31 34 -27
rect 27 -39 31 -31
rect 47 -39 51 -22
rect 0 -47 4 -43
rect -1 -51 3 -47
rect 7 -51 11 -47
rect 15 -51 19 -47
rect 23 -51 27 -47
rect 31 -51 35 -47
rect 39 -51 43 -43
rect 47 -51 52 -47
<< ntransistor >>
rect 5 -43 7 -39
rect 15 -43 17 -39
rect 24 -43 26 -39
rect 44 -43 46 -39
<< ptransistor >>
rect 5 0 7 24
rect 15 0 17 24
rect 24 0 26 24
rect 44 0 46 24
<< polycontact >>
rect 1 -14 5 -10
rect 11 -22 15 -18
rect 20 -30 24 -26
rect 40 -22 44 -18
<< ndcontact >>
rect 0 -43 4 -39
rect 27 -43 31 -39
rect 39 -43 43 -39
rect 47 -43 51 -39
<< pdcontact >>
rect 0 0 4 24
rect 9 0 13 24
rect 19 0 23 24
rect 27 0 31 24
rect 39 0 43 24
rect 47 0 51 24
<< psubstratepcontact >>
rect -5 -51 -1 -47
rect 3 -51 7 -47
rect 11 -51 15 -47
rect 19 -51 23 -47
rect 27 -51 31 -47
rect 35 -51 39 -47
rect 43 -51 47 -47
rect 52 -51 56 -47
<< nsubstratencontact >>
rect -5 28 -1 32
rect 3 28 7 32
rect 11 28 15 32
rect 19 28 23 32
rect 27 28 31 32
rect 35 28 39 32
rect 43 28 47 32
rect 52 28 56 32
<< labels >>
rlabel metal1 -5 -14 -1 -10 0 a
rlabel metal1 -5 -22 -1 -18 0 b
rlabel metal1 -5 -30 -1 -26 0 c
rlabel metal1 52 -22 56 -18 0 out
rlabel nsubstratencontact 52 28 56 32 0 vdd
rlabel psubstratepcontact 52 -51 56 -47 0 gnd
<< end >>
