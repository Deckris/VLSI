* SPICE3 file created from homework1_1.ext - technology: scmos

.option scale=0.01u

M1001 out in Vdd 0 CMOSN w=300 l=200
*+  ad=19000 pd=1800 as=19000 ps=1800
M1002 out2 in out 0 CMOSN w=300 l=200
*+  ad=19000 pd=1800 as=19000 ps=1800
M1003 out3 out2 Vdd 0 CMOSN w=300 l=200
*+  ad=19000 pd=1800 as=19000 ps=1800

.include tsmc025.sp
.param supply = 2.5

*c2 out 0 1pf
*C1 out2 0 1pF

Vdd vdd 0 DC 2.5

Vin in 0 DC 2.5

.tran 10p 1000ns

.control
	run
	quit
	*plot Vgs2
.endc

.end 
