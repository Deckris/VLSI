magic
tech scmos
timestamp 1639397274
<< nwell >>
rect -30 14 6 26
<< polysilicon >>
rect -25 18 -23 30
rect -17 18 -15 30
rect -9 18 -7 30
rect -1 18 1 30
rect -25 -1 -23 15
rect -17 -1 -15 15
rect -9 -1 -7 15
rect -1 -1 1 15
rect -25 -8 -23 -4
rect -17 -8 -15 -4
rect -9 -8 -7 -4
rect -1 -8 1 -4
<< ndiffusion >>
rect -26 -4 -25 -1
rect -23 -4 -22 -1
rect -18 -4 -17 -1
rect -15 -4 -14 -1
rect -10 -4 -9 -1
rect -7 -4 -6 -1
rect -2 -4 -1 -1
rect 1 -4 2 -1
<< pdiffusion >>
rect -26 15 -25 18
rect -23 15 -17 18
rect -15 15 -9 18
rect -7 15 -6 18
rect -2 15 -1 18
rect 1 15 2 18
<< metal1 >>
rect -26 22 2 26
rect -30 18 -26 22
rect 2 18 6 22
rect -6 11 -2 14
rect -6 8 6 11
rect -22 2 -2 5
rect -22 -1 -18 2
rect -6 -1 -2 2
rect 2 -1 6 8
rect -30 -9 -26 -5
rect -14 -9 -10 -5
rect -26 -13 -14 -9
<< ntransistor >>
rect -25 -4 -23 -1
rect -17 -4 -15 -1
rect -9 -4 -7 -1
rect -1 -4 1 -1
<< ptransistor >>
rect -25 15 -23 18
rect -17 15 -15 18
rect -9 15 -7 18
rect -1 15 1 18
<< polycontact >>
rect -26 30 -22 34
rect -18 30 -14 34
rect -10 30 -6 34
rect -2 30 2 34
<< ndcontact >>
rect -30 -5 -26 -1
rect -22 -5 -18 -1
rect -14 -5 -10 -1
rect -6 -5 -2 -1
rect 2 -5 6 -1
<< pdcontact >>
rect -30 14 -26 18
rect -6 14 -2 18
rect 2 14 6 18
<< psubstratepcontact >>
rect -30 -13 -26 -9
rect -14 -13 -10 -9
<< nsubstratencontact >>
rect -30 22 -26 26
rect 2 22 6 26
<< labels >>
rlabel polycontact -26 30 -22 34 0 A
rlabel polycontact -2 30 2 34 0 D
rlabel space 2 8 6 12 0 OUT
rlabel metal1 -26 -13 -14 -9 0 gnd
rlabel nwell -30 22 6 26 0 vdd
rlabel metal1 1 8 6 11 0 out
rlabel polycontact -18 30 -14 34 0 C
<< end >>
