magic
tech scmos
timestamp 1635696861
<< nwell >>
rect -11 11 3 21
<< polysilicon >>
rect -5 16 -3 18
rect -5 -1 -3 13
rect -5 -6 -3 -4
<< ndiffusion >>
rect -6 -4 -5 -1
rect -3 -4 -2 -1
<< pdiffusion >>
rect -6 13 -5 16
rect -3 13 -2 16
<< metal1 >>
rect -6 22 -2 26
rect -10 16 -6 22
rect -2 9 2 12
rect -2 5 6 9
rect -2 3 4 5
rect -2 0 2 3
rect -10 -8 -6 -4
rect -6 -12 -2 -8
<< ntransistor >>
rect -5 -4 -3 -1
<< ptransistor >>
rect -5 13 -3 16
<< polycontact >>
rect -9 3 -5 7
<< ndcontact >>
rect -10 -4 -6 0
rect -2 -4 2 0
<< pdcontact >>
rect -10 12 -6 16
rect -2 12 2 16
<< psubstratepcontact >>
rect -10 -12 -6 -8
rect -2 -12 2 -8
<< nsubstratencontact >>
rect -10 22 -6 26
rect -2 22 2 26
<< labels >>
rlabel metal1 -6 -12 -2 -8 1 gnd
rlabel metal1 -2 3 2 7 7 out
rlabel polycontact -9 3 -5 7 3 in
rlabel metal1 -6 22 -2 26 5 vdd
<< end >>
